`timescale 1ns / 1ps

module CPU_C_tb;

reg clk;
wire [31:0] PC;

CPU_C test( .clk(clk) , .PC(PC));

initial 
    begin
        clk = 1'b0;
        #20;
        forever #20 clk = ~clk;
    end

initial 
    begin
        #1000; $finish;
    end
    
endmodule
